module Instruction_cache (
    input [31:0] instruction_in,
    output [31:0] instruction_out
);
    
    assign instruction_out = instruction_in;
endmodule