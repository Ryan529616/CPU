�Ii2�*�� É"�t��kd�u� ���]yX�qq=�[�K��5)�Y�M�ש�}�f���#���w9��*n̲���(�,1 ��@u}�F`z~��K���SI;���y!j�1M`��<��Y@4����WK�i��SL�ׅM��^��|� $*��D%�&���~ϕ5�I�[t?c(���tD�+�!������U��X�ix��|������b�y��� 0!�؟{���C[��PZ�U��x5��|ά�h��P�!������At��hL���C�ᮗ˼^��t�)C>��(1ŕ���W�eN��|�\�.�j=z��U��S�����e�|���D��>o��Ӯ�_��)�W����~[� Y6G1lڄ9,�d�Qq���H� � (�s�}��nu����y�I	ђ#f9��]z�|4ib��i�K��	��M{�pu�xf�ߡ��|��d31҇��sH%�Or��烔��+Ct7 ����G{˫`]��9�3���K�����w�Чs�y.1)��!��H?�W��#e?@�ɹ�cjȞ�q���P���������&�AV暑���s���wvz�:#��w߀�����I$j��_({L��i�F�:��R�w�% �u�_f��i����ix�`K��Ņ5g4#LK�\/���"'�O���ɚ����1�+Y���R7�c ,.L�E�}��y^k±,Er/��kO04o@ Ө����9�) �M�U4�4rW���!t�,ARR*��{5�h�� ����K�������VK��m|�����:�)	�?����EjTG������#��{��p��\�Y�5�4٦�%�h�:&p�wM~0�"�Eٟ�K9����-�:bC:��_u��5i��J�1V!8�S�c���wٹ�����V>��n����4!'ydQ$s�0+� ���Xv�O8Y���<B�zf���~��(k���D��Rq�a17��Y����B'#w��Y2��:������ڲ�&�����'c��G�̲Z���kV)l��w{V��I���+ظ�Q~�����p�9i  �#���o�G<s��<�)`������ܠa*Ma���hQ�G��?��I��9w��QCR������G�b��-EY�7'w�.��`ͅ}%-�v�>q�+����.�ȇ�!��.s���ۓ
�t����z�ګ�*��m��^�u�5)nz�	,�Yk�=�
��Y��"��JY� $s��*C��>���/خ�yk��>��L�W���ġw]Oቭ�$�4�X���Q� �lM�+�!�8f�5}�k\o�\Os]����ۜK��S����dKz`w��9c�s$��F�C����!��+�cY����g���`�JŐ����ʗ�^oH��#n�w��b&�1>Q�3��u�A�r���!����6�
A�ى��u����EX[����\S�yaB�����NR��v���IS0��¨H�'B��1x� kʈ>gr����hӗ5*U2��w[�m�/�@N�%�ۚ�^�;4�%���;�h"���	(�8;=���h�bcE�$���q�jdw�[F���)��~wn3�~�C���
���Ē0!�y+6>PW�%��O���)��AD���I����&<t`�_T�qΆ�����.�'�i�����}�� pɕyh�|���k�����N�9X0�w3=2�χ[�i��|v\�ӧ��R�Y~���Ɲ��-f��j�w�PC�-ULN�"үe��:���mܕ�#�+���v��0y�����{r�)�����Y�^�~gS�y���Q��NXF�]'��Ew����Tc���T��n-��&$�X����_��A&S!���g�r��N�SI|��F�@��O����ũ