�Ii2�*�� É"�t��na�p�%���X��q�K�X�[	y�q=��Q�+��$�@��Ъ^C�N_:��.旌��F�R�S ��p��~v4�͢N=�#.!�bx��bv"��=��q�+�l�#X�S�u��ژ�N��NWk�Mee�����m�U���ј��8۫Kq�Y�j��|t�44��V�]vq�]\VXL�^|}�lP�F�!bY��ڵ&卄6��`����?xɥ*1I'��
>�D��K��B����f�1<���jT���rB�q���X�I�� ��;�ϪL1�L�k�m2נA�I>F���]�+N�
��<s]���κj�4�6`{�8�$�_��`��<r�ԏ��&����[F@j)��sJU�j��{���9���2р��X������3
��G�RN��似��E �6h�;�,lqxv���1���������	*�J�G�.����"����v�3������4[�ɗ,�8������Dw��Ĳ{R5]�g��תR������G}S	�	L�ŧЕ������}��E���ۓ6���Z'K�\����-$���e�b<��L ��NՍj�SKu`�:4�L�z·�m+��yǁ���S���C��O���/Ǒ�5�#e�B�͈����˅I��V� �C6�����CA~���%�,Z�
A�����_o���Z�1W�]���M98LQx?0�/��+����(`K�#ۅ��8��{u%P�� A�� ����ǭ�gF���im�V	t�+�?R�~��b�2w&���rT>�'�P���2&������t@���ԑ�.Xto����@�I�@p�*�G��������Wtb7�b��
C�7��?{_�F�`�;a��}�E6B	.�PO��-��&��:�in�q�a����ɫ�_5�
?Q:<e# H��E��L���䘴fY W��3P7H(��.-�R
_M�� u�W��-����=��Jx�>��6-3��ʂ���01��*��~�e׳����ԏJ�08.n!��e�3D� E<��ك�'Ӈ[BY���!�<��r��`Όʼ|�lPngF�Bw�Ys�'��q	�� 05(!�]sh<Nq_22�&��!���`�B�e$ώb��Xs`�^n��m�)�]���wvg��;��c��S��{�@���ʻcr[�b��"�8�ڨ����t+g[�"����A!�E.�K��`�z��=��H�Y���<L�m�U������+>�	$�jeשQC�FOk����,�l�V����z�yi�î�"��[�Lu�'�KHV�d���ES��J�b���Q�]�}��J֞�!�f�(�9��I٠�S�0a$��rG��y�On K���W�H����[S���i��l�� �B��g�\7�����QK������pM*	�$�yu�u��>sh:�{s:���ϭ��gd��G�J ��d��ej�ke�$2�V~�r¨�4Ur>�T��ќ���t�C·��}��%�"��e;Yu��P^Ԇy_�c�d��#��]����OIUˏ�h(T��ᤷ}�U��k���S5�`������tZ�S4+5a�{nۨ�Fn����@J	-S3��Y�S�+��CX�_Be�%l��$�D�?���P^�!��	�@fZ٪˝��f�a�]Eo�J �D>j"uC�a3�WX���X��܆�����@r�t�M�	@a#�N�����%�S�����mD,
"����8u14��`���K̴a�k��[�V��$fx�k�&7>7_i2\j`A��4�CV�0L.X�)ٖ�i"oX��>�CX���4����PbUTh��uxN���Ā����C�;�Qѳ�ѿcÄ��9��Q�G�/�h���o�L�wSP _����T��E5"���#�����@�{nc�TN~"��O>R��fPl�4q��r<��}�1+j֍���~Za1�,�]��,D0�c��oLp�����b[*1�g���H`:4gw�3��XXX_-���ˈ�����"�Un���ʬun�k0��=il
�h�*�!���U�v���v�ܥ�6���Ļ�Þ�l�?.�؝��ׁ����]�|�Ă���8��{LL� )�h/wv94X;~��O%=�+='�m�`G���a�HF�|뻬�ꉖ�!5��� {�p�zre��]���?Xh~��7n8�V�g5��AiV����D�汩f��W�c��[0�,�ů���2Fab�i�Ѻ�5)V����_�Y^,������OQn�r͐s�����~�>z��k���D�(�=T�7���6���>O�7���[��$̇�,��ߖ�r����ԑN�V�ϕO}�Pq�8����vg�v��n�p��~��̱����K�1(D��,�Dr�?~:�J��)V�d�|Tf�G�3�B�����*��>p�(��ػ��w�⻕��͟�7��Dj☻'$'X���7�ZάN�-oM���y\U��{�bD���$��h��Ε�+�ߞȗ�K�-A�ƞ��MZ#��r{���|Q�)����t6o�d��~iE�Fєi�Xl���`�Id�_�YĪ?�~O�\u��%O�|�j6��`�Ѣ��@���k���wy�NQ(�6�1Y`���b��,�>�~,�7��2!�R�k2�I׀$�o��+���t造�~Z����E��O*~_�<�3��uV�v�=��6�A"'��݉l�%�JJ�(*l%��k��E͝�8�,,�G����L�b�p� �~�Eov�^-i��jd�ڈ��`��}��9e��^����ۢ�A��ǎiJ������W�Z���̃z �f����SiXJ������i��`<�~ <vn
��,C⼜N�V�����TN�����S�G�<1��?f�#!��#˵o@���jБ���dR֘�o�� �*km��g:�O�[�z,V�*>���B�U�BMcT�oA=<s~����ei0l|���@�2m�RU�Am+���i5�]�?M��rs���m��r����+=�a4�"�k�����S���d��^��r�٤iQ�L1�\-��^G���5�3??,pdJ'4�b$�HW[����<�����t�)`=MK�˝���(of��8;<�$\�¬'fs�Vp���ٗ��gi��S���Ѥ��q�;�0�J�K�C�e��&����x"�(Ս�+җE&X�Z��$:Qt4/ ����@c3Ǎb���K��i�RZ�T�� >������wkbsEƹ���/>
�2��G��\��7�����H��~E�;ݓ�$���:x˓�3�y���4�e2��
k����d�K�/��L3)J�<�{��2��νK��/�6ry�u~�z�^���J�rh���ICI�@#M���ts�ܻ��yҀ]o�� ]�8@�g~��7�������]��Q-l�a�{��ps�?nC$Xd5� �Z����;v��ȄtM��ov1>$��+�'=�w\"�����ygt�e�HpG���%5����$�*1g��Ǿ�m�V���_�����ں��u�b���S�fG�
5HR8��.[÷y~kw�x��NϿ���4D/�:��]
����D�V/�ׄ�媞��G���2d�_��ٚ�ȣ$�\�%o�B?��XpjCb�I��іO`�7�����	$�@A�A���j����E�G�́˸�ˍ�UU*B���7!�ܵ����=:4�HB��ހ�g��<i��}���#8��~9m-�[,k@���5�%�SS	�k��`�􀳣�ߖT�n��Ѽ�n ��t��\I�2umgh����kL��p+pm�+Rw�k�HD}�L�[p���̿Z���O�2.`YcX(����%�\訪%K�(��v�� �S#�G(ĺ5v��'�^mH4	�� ��7�"�C ��>I��sWp췰Bq2 ��L��*�5�4-�WŉX� <�����*k���ҩ��˼L�>r����� �xժP�o:P7��!�s�������$�����v�~96�f�f�k�$(dU^_�>5_L��|T'y�?h���h��d�"WU���l��v�s1ЃgK̈́X�>�����X���G�U0;�r�#  ���y���߅q�J��ܤYm�1!t�E���/2�^�H7�����!����3�W�t����9�h>Q��(;�\\����J��������D-�I�N.��}����L{9)��׎p��PN�jE̞�Z��P]��r�`/+]> ������,J���w����T�l��a%��$N�lP �q��ՅΥfxn�ɚs�ƾ&-�|x�x�,��;w ����I���F�<L�IFyF�ON�V!���fX6�uZ�,6��>Pj�kW�w�T���NƐ�;$��x�@�s�y���L��DQ�E]�2�؇��8���^�2�])D��@�������n��!���('��B��m��� �wC�0�\�z~�}�<�=dy(�'qcf�T��Iys�;R�Ũ�P>��������p��*�b��E�/S�eo���a���|��%ό?#��`�
���l�Vl���L%Ep.0%3�E6>�`�Y�Lf��8���<��n�u�II^�ˌ͉�ҟ���X�O A�@*sWU�-�v���O�bք񂁙X@}�ղ�n_	�x�Y��8E��g��
+�(^�E�1߲#oWTZ� ��N�K=�%�/1�Ũ�"��N���n�N�F�����әPU��z'�����*8��ψ�G������Dg���+J�?'g�̈́���"^ȓgHȫ�@<��Xbؼ@�ZF�A�J��z�a��f�Z؆Y��~nz����AT��Lp�=�E��Ђ�w���;�=�C"�?/�<wo�NH���)�^�(u�|͐�U5E�sʥʊČ�,���~5�ODo��a��l;���:�:�*�� �<.ϽF壞l����
��G��N�@VLJg�t��� J�OOj��I(����$^ė>��㋚X���r��F`���bǐ��$i�*��C���(��j����E�n��=��C�Y߭<ր~U��ˆC�z��:8��/0��4��3zi�� �??�gb9*���3���(���-�0͏ΰ빀4{
��
{��	#������Dd0�� �������m�~~�����������j�`k��HԱ5�%d$/?�h݊h�Sy^G��Y�A��:#��e%��#S�kA6g��d��`yf.|M�� ���L�I�Rf>(����c�!�K�S�����6����\q�B^�����_-�����ᕊ\�m�VX��ٻ���/�t��;�;�^0�#��[L�q,���� �-S�l�i�M�-�j��-YH��p�EX�"A�#���`���,G�s\���]���9���Hhm3���߯c�ky�B��@l�`�a��N�T��]ˌA�_(k�߉���m���K-m΀���9{@�DH��	]�\�M��]�'��;1��0�<`��ٔsV�Fˉ�J&��?������=H�N[a����B�q�3��Ք� 4�+�w9F��+Z���1����$��뺌���״,�g�=T<~]I0�ϖyZxݰ\璅�r
,�,s %BM�y� �"�ZB�9`g�i�&��;%I�F�,���)A�f �9�\�2+��pJ$G�rn��<[�Qt�}�X��$������CTϱ�W�M�k�[�j�T�E���!H�y8M�
��َ
c�#���o�˅ӑ�8>"?��/0��7���U]mi1`���6�6�(^��/�nvE\���1[�I��Җ{�����/뿝I��i(�R�^��e����b����];c�q���;G�n�q�-N�Fc��B���=�cB�������� pgͨ6v��9C���׷���LK����D��d� ��]&�"ݟ%�GFjYֻ�zV1~s�4�ds���&bXv�H�B�J�}M=�D�����r6>
kH
������d��?�*���L���e5��S�TT��;%%��[R��e������l
;�"�θ�f禽�kX��#�+�L8Z�@������A���G'U��x�V����8���?�5�2f(���y���x	��dU�q�c��)nYX:�V�S�7��*�X���5��Yb�4��݇�)��'�{a�dK�BPE{�)�{��)kdO�;p$%�í� 0S�*6�*v���iV|KX����l�����Q�RnoE\R�Ň���(�R�v_��w���99�;f�!ML !��E(��G���9�_�#��.l'���Q2��p�R݁��H����]u��4��hee���ѻ�W]IG[@֚�J�bZ�����-������W�&���<$ħ̃��SM��R�8��HLg��,�{���ck��ȥ��n��4ہ���U�����3l%ϛ�)�X� ��ŜA?�+�h_��V6��,�gY yKq)z(�]��/�3����%�iRs�M|ǽ y_�0eAѲ��X��PƬ��.dsX�
8}ٱS����h�15�ٹy� �g�K������>BZfM|X����Dܭ����q�i�plE��.˟��D�*.(B�'�<ET,���%�-�>j8>fe!XL[�:��:�(���qŠH	4C՚OU�YW~�	Dx*i_��7�e�
;����
�i��k(��m�hX9v�������$���M�n?���Tu�o��O���_H�-t0��r]Qp}��[�j�1|#-����-���qU��p��nb�P�� 
��LT���S�c>���E#���@����Y4������:1�����ןm�q��٩�8��آ��W!;���-o����p����O���{�����r��\ȝ�8+��gY��7;����^ťF�F0��ǳCد���@�gn�*��8P�\�� 	�٧$�!�G�/�X�&_2�حڠ����s�,� �}�)�h��E��#��N�R�spn�x���)�h���H�7���W
�?�������o�)�4]kn�M�McY�~�v��r���H�qQz�w�;��f$ٛ�c�����r.���Ζ@wFQ<^ߣ�w�Hv+*�=;ڛ|�����Vx�J��EC<�.�����!1ͣ]�{�_�hM觔��E��M�Am���{�c�d�IY)o���,rՁ+�K���"ylB5C��:9�E����:m�)؈*U��f�Z;2����5�m̆��=��Ƈ���uEk�#����<�n���yr�zfXq��{�'+���c$�	a�.�>:~ߪ��y5�%���6�t݆���ep6�ꅈ��%��s�	�׸�/W��9�y<�%����c�J�Y�������t�N-�l�d�S'q�w�<�1�Ev�Z]��z��(M��{6_8ҷ�4��ҥ0a@�������;z��r���Y^l
#��0�$s�����ޛ�V!ϙ�N��M��݇d��Q�^] ټ� 1(�]�ŀC���r��_F3y���	WNy@ռ�.�� �x���L7F�֠)6���M#kʮ�꣒���W�w��Lш�y�)�w� �Q��l"j3Z7Y�*����8�wS�y��S@8�>)-G�0�9�Ou5���eY�oh���B�cf���^��;��!GKx�!�$��p�	9�H��o��I䶑�E�[�A.Fn�D��UPZ���wP����2+�˿��:������e]��:'H��U��=D��\X7w��\�O3��c��n��	aM�k���p®� ���F{�=})6_�L=���~��x�LK2��}UMr-��h�+�+#Z ������oA�c���Q-f�3�!��A�]+�j�i��k�$X��>�ѬO�A�cwSM�T�po-�,���XqvƮ�!Q٠&�#mFW����udSl��usgu��Hj��kɚTῥ���bd�j���Q{��Y.x[?�S>A޶���]E��wZ���Ϥ��ɠ�J/x��V�|qߍd����si>h��ѻ��R���M��%�[�(y��mOu�7�l��*��ɔ����1�;:^j.��5J��!�)�����B�R|]0.!%{V(��ç>Pa1��T%�S�v�+Ҳ�eSfQ��%a�{��?�N�}�|���sp��T�Ɯ���/(FZ[G�L��������b.��^��b�,�F@4>��N~��.@nV���c�*�$o�C���)��}3�Q���`�>ʧ0lc�S�S�ϭ���UZ}�1ȘǓ��y�4adp�Wd�@�<,G,�ë���fC�R��;~-�W��\�0�Y��Tq<���`����F��-�o\}uPU�$���ŭK�*�v�����Xt��_S�,�i~�]�{�4�8�K��@�,^Pz��L:���ݦw"������z��[��Μ�����f��gQ�s�g��l�j�H)Q8�E_��e]�9��#x]�]Y�M�]P�L(�����^���
7�Թ����x9�;�����C��}�X穾zY�]�����h8���XR-���`�¥ۋ�.�\��&�[T���*]��|���!�����I	����Է�����h0D��Fifo�DK+ ��Ы+۽�#WTau�ύ�W��0��#r+�5޿����l��C�F�����WB��yC�����a&(	���7^jr'��Kњ�H��N�%�c�&���	��mO���s/�f�H��f�<�H:L�[@��z.?�A3�A[��,?["S�mL8$�d
�0�_��O�����:%��n��������L-$:&�G�y�|�����kо�y�iS�'��̾��-�=)�ę-C��#�bE�\�~V2_��<b��'K�m�@"x�$6�6�N�������jU�Ֆ�S��8R�@���cy5\U��������1#��y��=TQJ� ".��-��M��Y{.,3:�b˱꒯j~��X�4�̃(x��3+Y���G���Pck���I��>4�T��r}e1ȩ� �jO�7̟!�G�W�n���M-�n=w_�J y?�=�v�;t�W����E�N�M��t�T<�l�ƹ��΅u*~"8kV|��?�<�N�mr��]��%F�ǖ��K�Lq���A�����Nm��8V+�h�X�U���+Ѩc�#D�M�ZG�}�d1��/j:�SN>�LI��!���s2MX�ً9g������j#U���F����e��іj�	[�y�@x'W����^�=��&�z�mL7&��\�1�Ŀ+Kl\Ҽ��cX�7����y~S������l��ec+k��ܴJq+k^��|��)��YQ����/����kM���OR�8����վ�Rk9�{<[��ɺ0��-93�@�-��	2�`�����ڋL�l�%��<�~N���7y�;��Ă�F����a8KXI��K���T\�f$_�&N����ݼe��$.�.��U.G �${^�c'�^��Q2�ˍ�|��q;�5��QC��Yv�= �w���Vb'�B���#����t*���o�v�V�2��m��~8��'��<=�?�,3d� gK����A ;d(]��ڃ�$����E��J�l��Pr�.�K����w$Ȋ5_�2H_���d�'@xc�z���%�D�Z���0�U ����"�3Tz������&�e��.�A��e���wl��Pu"�Z�I���ݵ��є?�ԘƂ�b)1�8��C'�"Wo�^�m�3.'�%{TK�Hr��@�ܱ<� Ϛ݉¤��LX����!��̥�A�����545�ED�b}]���G왟t�Q��˃U�C��b�l�˾�{ 